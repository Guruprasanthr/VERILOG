module pe (
    input  [3:0] d,
    output [1:0] y
);
    assign y[0] = d[3] | ((~d[2]) & d[1]);
    assign y[1] = d[3] | d[2];
endmodule
